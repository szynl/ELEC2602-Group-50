module binary_to_7Seg2(binary, sevenSeg);

	input[3:0] binary;
	output reg[6:0]  sevenSeg;
	
	output[6:0]  sevenSeg;
	assign sevenSeg[0] = ...;
	assign sevenSeg[1] = ...;
	...
	
	assign sevenSeg[6] = ...;
 
endmodule
