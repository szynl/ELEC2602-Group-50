module instantiate_lab4_part2(SW,LEDR);
 
	input[9:0] SW ;
	output [9:0] LEDR;

	// instantiate and connect master_slave
	
endmodule